module ram_controller(



);



endmodule