module dumpvars();

initial begin
    $dumpvars(0, bits_testbench);
  end


endmodule